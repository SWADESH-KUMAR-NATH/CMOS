*Divider CKT
Vbat  vin   0     DC 5
R1    vin   Vout  1k
R2    vout  0     1k

.control
tran 0.1u 1u
.endc

.end

